magic
tech sky130A
magscale 1 2
timestamp 1679616029
<< error_p >>
rect 19 481 77 487
rect 19 447 31 481
rect 19 441 77 447
rect -77 -447 -19 -441
rect -77 -481 -65 -447
rect -77 -487 -19 -481
<< nwell >>
rect -65 462 161 500
rect -161 -462 161 462
rect -161 -500 65 -462
<< pmos >>
rect -63 -400 -33 400
rect 33 -400 63 400
<< pdiff >>
rect -125 388 -63 400
rect -125 -388 -113 388
rect -79 -388 -63 388
rect -125 -400 -63 -388
rect -33 388 33 400
rect -33 -388 -17 388
rect 17 -388 33 388
rect -33 -400 33 -388
rect 63 388 125 400
rect 63 -388 79 388
rect 113 -388 125 388
rect 63 -400 125 -388
<< pdiffc >>
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
<< poly >>
rect 15 481 81 497
rect 15 447 31 481
rect 65 447 81 481
rect 15 431 81 447
rect -63 400 -33 426
rect 33 400 63 431
rect -63 -431 -33 -400
rect 33 -426 63 -400
rect -81 -447 -15 -431
rect -81 -481 -65 -447
rect -31 -481 -15 -447
rect -81 -497 -15 -481
<< polycont >>
rect 31 447 65 481
rect -65 -481 -31 -447
<< locali >>
rect 15 447 31 481
rect 65 447 81 481
rect -113 388 -79 404
rect -113 -404 -79 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 79 388 113 404
rect 79 -404 113 -388
rect -81 -481 -65 -447
rect -31 -481 -15 -447
<< viali >>
rect 31 447 65 481
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
rect -65 -481 -31 -447
<< metal1 >>
rect 19 481 77 487
rect 19 447 31 481
rect 65 447 77 481
rect 19 441 77 447
rect -119 388 -73 400
rect -119 -388 -113 388
rect -79 -388 -73 388
rect -119 -400 -73 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 73 388 119 400
rect 73 -388 79 388
rect 113 -388 119 388
rect 73 -400 119 -388
rect -77 -447 -19 -441
rect -77 -481 -65 -447
rect -31 -481 -19 -447
rect -77 -487 -19 -481
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.0 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
