magic
tech sky130A
magscale 1 2
timestamp 1679616566
<< error_s >>
rect 1695 1254 1753 1260
rect 1695 1220 1707 1254
rect 1695 1214 1753 1220
rect 180 881 238 887
rect 372 881 430 887
rect 180 847 192 881
rect 372 847 384 881
rect 180 841 238 847
rect 372 841 430 847
rect 492 832 514 900
rect 926 851 984 857
rect 1118 851 1176 857
rect 84 653 142 659
rect 276 653 334 659
rect 84 619 96 653
rect 276 619 288 653
rect 746 638 768 832
rect 926 817 938 851
rect 1118 817 1130 851
rect 926 811 984 817
rect 1118 811 1176 817
rect 830 623 888 629
rect 1022 623 1080 629
rect 84 613 142 619
rect 276 613 334 619
rect 830 589 842 623
rect 1022 589 1034 623
rect 830 583 888 589
rect 1022 583 1080 589
rect 1599 326 1657 332
rect 1599 292 1611 326
rect 1599 286 1657 292
rect 971 279 1029 285
rect 971 245 983 279
rect 971 239 1029 245
rect 450 232 508 238
rect 450 198 462 232
rect 450 192 508 198
rect 971 -231 1029 -225
rect 971 -265 983 -231
rect 971 -271 1029 -265
rect 450 -278 508 -272
rect 450 -312 462 -278
rect 450 -318 508 -312
rect 881 -635 939 -629
rect 881 -669 893 -635
rect 1546 -656 1604 -650
rect 881 -675 939 -669
rect 327 -683 385 -677
rect 327 -717 339 -683
rect 1546 -690 1558 -656
rect 1546 -696 1604 -690
rect 327 -723 385 -717
rect 785 -945 843 -939
rect 785 -979 797 -945
rect 1450 -966 1508 -960
rect 785 -985 843 -979
rect 231 -993 289 -987
rect 231 -1027 243 -993
rect 1450 -1000 1462 -966
rect 1450 -1006 1508 -1000
rect 231 -1033 289 -1027
use sky130_fd_pr__nfet_01v8_J2SMEF  XM2
timestamp 1679616253
transform 1 0 1000 0 1 7
box -73 -288 73 288
use sky130_fd_pr__pfet_01v8_XJKEBL  XM3
timestamp 1679615849
transform 1 0 1003 0 1 720
box -257 -150 257 150
use sky130_fd_pr__pfet_01v8_XGEZDL  XM4
timestamp 1679616029
transform 1 0 1676 0 1 773
box -161 -500 161 500
use sky130_fd_pr__nfet_01v8_PL7QEV  XM7
timestamp 1679616029
transform 1 0 1527 0 1 -828
box -125 -188 125 188
use sky130_fd_pr__nfet_01v8_PL7QEV  XM8
timestamp 1679616029
transform 1 0 862 0 1 -807
box -125 -188 125 188
use sky130_fd_pr__nfet_01v8_J2SMEF  sky130_fd_pr__nfet_01v8_J2SMEF_0
timestamp 1679616253
transform 1 0 479 0 1 -40
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PL7QEV  sky130_fd_pr__nfet_01v8_PL7QEV_0
timestamp 1679616029
transform 1 0 308 0 1 -855
box -125 -188 125 188
use sky130_fd_pr__pfet_01v8_XJKEBL  sky130_fd_pr__pfet_01v8_XJKEBL_0
timestamp 1679615849
transform 1 0 257 0 1 750
box -257 -150 257 150
<< end >>
