magic
tech sky130A
magscale 1 2
timestamp 1680540636
<< nwell >>
rect -257 -150 257 150
<< pmos >>
rect -159 -50 -129 50
rect -63 -50 -33 50
rect 33 -50 63 50
rect 129 -50 159 50
<< pdiff >>
rect -221 38 -159 50
rect -221 -38 -209 38
rect -175 -38 -159 38
rect -221 -50 -159 -38
rect -129 38 -63 50
rect -129 -38 -113 38
rect -79 -38 -63 38
rect -129 -50 -63 -38
rect -33 38 33 50
rect -33 -38 -17 38
rect 17 -38 33 38
rect -33 -50 33 -38
rect 63 38 129 50
rect 63 -38 79 38
rect 113 -38 129 38
rect 63 -50 129 -38
rect 159 38 221 50
rect 159 -38 175 38
rect 209 -38 221 38
rect 159 -50 221 -38
<< pdiffc >>
rect -209 -38 -175 38
rect -113 -38 -79 38
rect -17 -38 17 38
rect 79 -38 113 38
rect 175 -38 209 38
<< poly >>
rect -159 50 -129 76
rect -63 50 -33 76
rect 33 50 63 76
rect 129 50 159 76
rect -159 -88 -129 -50
rect -63 -88 -33 -50
rect 33 -88 63 -50
rect 129 -86 159 -50
rect 129 -88 225 -86
rect -159 -97 225 -88
rect -159 -118 175 -97
rect 159 -131 175 -118
rect 209 -131 225 -97
rect 159 -142 225 -131
<< polycont >>
rect 175 -131 209 -97
<< locali >>
rect -209 92 209 126
rect -209 38 -175 92
rect -209 -54 -175 -38
rect -113 38 -79 54
rect -113 -94 -79 -38
rect -17 38 17 92
rect -17 -54 17 -38
rect 79 38 113 54
rect 79 -94 113 -38
rect 175 38 209 92
rect 175 -54 209 -38
rect -113 -128 113 -94
rect 159 -131 175 -97
rect 209 -131 225 -97
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
