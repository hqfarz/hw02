magic
tech sky130A
magscale 1 2
timestamp 1679616029
<< error_p >>
rect 19 172 77 178
rect 19 138 31 172
rect 19 132 77 138
rect -77 -138 -19 -132
rect -77 -172 -65 -138
rect -77 -178 -19 -172
<< nmos >>
rect -63 -100 -33 100
rect 33 -100 63 100
<< ndiff >>
rect -125 88 -63 100
rect -125 -88 -113 88
rect -79 -88 -63 88
rect -125 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 125 100
rect 63 -88 79 88
rect 113 -88 125 88
rect 63 -100 125 -88
<< ndiffc >>
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
<< poly >>
rect 15 172 81 188
rect 15 138 31 172
rect 65 138 81 172
rect -63 100 -33 126
rect 15 122 81 138
rect 33 100 63 122
rect -63 -122 -33 -100
rect -81 -138 -15 -122
rect 33 -126 63 -100
rect -81 -172 -65 -138
rect -31 -172 -15 -138
rect -81 -188 -15 -172
<< polycont >>
rect 31 138 65 172
rect -65 -172 -31 -138
<< locali >>
rect 15 138 31 172
rect 65 138 81 172
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect -81 -172 -65 -138
rect -31 -172 -15 -138
<< viali >>
rect 31 138 65 172
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect -65 -172 -31 -138
<< metal1 >>
rect 19 172 77 178
rect 19 138 31 172
rect 65 138 77 172
rect 19 132 77 138
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect -77 -138 -19 -132
rect -77 -172 -65 -138
rect -31 -172 -19 -138
rect -77 -178 -19 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
