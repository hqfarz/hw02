magic
tech sky130A
magscale 1 2
timestamp 1680477288
<< nwell >>
rect -161 -500 161 500
<< pmos >>
rect -63 -400 -33 400
rect 33 -400 63 400
<< pdiff >>
rect -125 388 -63 400
rect -125 -388 -113 388
rect -79 -388 -63 388
rect -125 -400 -63 -388
rect -33 388 33 400
rect -33 -388 -17 388
rect 17 -388 33 388
rect -33 -400 33 -388
rect 63 388 125 400
rect 63 -388 79 388
rect 113 -388 125 388
rect 63 -400 125 -388
<< pdiffc >>
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
<< poly >>
rect -63 400 -33 426
rect 33 400 63 426
rect -63 -431 -33 -400
rect -118 -438 -33 -431
rect 33 -438 63 -400
rect -118 -447 63 -438
rect -118 -481 -102 -447
rect -68 -468 63 -447
rect -68 -481 -52 -468
rect -118 -497 -52 -481
<< polycont >>
rect -102 -481 -68 -447
<< locali >>
rect -113 442 113 476
rect -113 388 -79 442
rect -113 -404 -79 -388
rect -17 388 17 404
rect -17 -446 17 -388
rect 79 388 113 442
rect 79 -404 113 -388
rect -118 -481 -102 -447
rect -68 -481 -52 -447
rect -17 -480 125 -446
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.0 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
