magic
tech sky130A
magscale 1 2
timestamp 1679615849
<< error_p >>
rect -77 131 -19 137
rect 115 131 173 137
rect -77 97 -65 131
rect 115 97 127 131
rect -77 91 -19 97
rect 115 91 173 97
rect -173 -97 -115 -91
rect 19 -97 77 -91
rect -173 -131 -161 -97
rect 19 -131 31 -97
rect -173 -137 -115 -131
rect 19 -137 77 -131
<< nwell >>
rect -161 112 257 150
rect -257 -112 257 112
rect -257 -150 161 -112
<< pmos >>
rect -159 -50 -129 50
rect -63 -50 -33 50
rect 33 -50 63 50
rect 129 -50 159 50
<< pdiff >>
rect -221 38 -159 50
rect -221 -38 -209 38
rect -175 -38 -159 38
rect -221 -50 -159 -38
rect -129 38 -63 50
rect -129 -38 -113 38
rect -79 -38 -63 38
rect -129 -50 -63 -38
rect -33 38 33 50
rect -33 -38 -17 38
rect 17 -38 33 38
rect -33 -50 33 -38
rect 63 38 129 50
rect 63 -38 79 38
rect 113 -38 129 38
rect 63 -50 129 -38
rect 159 38 221 50
rect 159 -38 175 38
rect 209 -38 221 38
rect 159 -50 221 -38
<< pdiffc >>
rect -209 -38 -175 38
rect -113 -38 -79 38
rect -17 -38 17 38
rect 79 -38 113 38
rect 175 -38 209 38
<< poly >>
rect -81 131 -15 147
rect -81 97 -65 131
rect -31 97 -15 131
rect -81 81 -15 97
rect 111 131 177 147
rect 111 97 127 131
rect 161 97 177 131
rect 111 81 177 97
rect -159 50 -129 76
rect -63 50 -33 81
rect 33 50 63 76
rect 129 50 159 81
rect -159 -81 -129 -50
rect -63 -76 -33 -50
rect 33 -81 63 -50
rect 129 -76 159 -50
rect -177 -97 -111 -81
rect -177 -131 -161 -97
rect -127 -131 -111 -97
rect -177 -147 -111 -131
rect 15 -97 81 -81
rect 15 -131 31 -97
rect 65 -131 81 -97
rect 15 -147 81 -131
<< polycont >>
rect -65 97 -31 131
rect 127 97 161 131
rect -161 -131 -127 -97
rect 31 -131 65 -97
<< locali >>
rect -81 97 -65 131
rect -31 97 -15 131
rect 111 97 127 131
rect 161 97 177 131
rect -209 38 -175 54
rect -209 -54 -175 -38
rect -113 38 -79 54
rect -113 -54 -79 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 79 38 113 54
rect 79 -54 113 -38
rect 175 38 209 54
rect 175 -54 209 -38
rect -177 -131 -161 -97
rect -127 -131 -111 -97
rect 15 -131 31 -97
rect 65 -131 81 -97
<< viali >>
rect -65 97 -31 131
rect 127 97 161 131
rect -209 -38 -175 38
rect -113 -38 -79 38
rect -17 -38 17 38
rect 79 -38 113 38
rect 175 -38 209 38
rect -161 -131 -127 -97
rect 31 -131 65 -97
<< metal1 >>
rect -77 131 -19 137
rect -77 97 -65 131
rect -31 97 -19 131
rect -77 91 -19 97
rect 115 131 173 137
rect 115 97 127 131
rect 161 97 173 131
rect 115 91 173 97
rect -215 38 -169 50
rect -215 -38 -209 38
rect -175 -38 -169 38
rect -215 -50 -169 -38
rect -119 38 -73 50
rect -119 -38 -113 38
rect -79 -38 -73 38
rect -119 -50 -73 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 73 38 119 50
rect 73 -38 79 38
rect 113 -38 119 38
rect 73 -50 119 -38
rect 169 38 215 50
rect 169 -38 175 38
rect 209 -38 215 38
rect 169 -50 215 -38
rect -173 -97 -115 -91
rect -173 -131 -161 -97
rect -127 -131 -115 -97
rect -173 -137 -115 -131
rect 19 -97 77 -91
rect 19 -131 31 -97
rect 65 -131 77 -97
rect 19 -137 77 -131
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
